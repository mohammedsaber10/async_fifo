class w_sequencer extends uvm_sequencer #(fifo_w_trans);
`uvm_component_utils(w_sequencer)

function new(string name, uvm_component parent);
super.new(name, parent);
endfunction


endclass
