module debug;
import uvm_pkg::*;
`include "../fifo_seq/fifo_w_trans.sv"
`include "../fifo_seq/fifo_r_trans.sv"
`include "../fifo_seq/fifo_w_seq.sv"
`include "../fifo_seq/fifo_r_seq.sv"



endmodule
